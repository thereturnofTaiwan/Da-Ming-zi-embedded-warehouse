module Flowing water lamp(
 );



endmodule
